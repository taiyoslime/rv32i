`timescale 1ns / 1ps

`include "define.vh"

module core(

    );
endmodule
