`timescale 1ns / 1ps

module fetch(

    );
endmodule
p